module arm (
    clk,
    reset,
    PC,
    Instr,
    MemWrite,
    ALUResult,
    WriteData,
    ReadData,
    DMSrc,
    ShftOp,
    Division,
    Multiplication,
    DivMode,
    NewInstr
);
    input wire clk;
    input wire reset;
    output wire [31:0] PC;
    input wire [31:0] Instr;
    output wire MemWrite;
    output wire [31:0] ALUResult;
    output wire [31:0] WriteData;
    input wire [31:0] ReadData;
    output wire DMSrc;
    output wire ShftOp;
    output wire Division;
    output wire Multiplication;
    output wire DivMode;
    input wire [3:0] NewInstr;

    wire [3:0] ALUFlags;
    wire RegWrite;
    wire ALUSrc;
    wire MemtoReg;
    wire PCSrc;
    wire [1:0] RegSrc;
    wire [1:0] ImmSrc;
    wire [2:0] ALUControl;

    controller controller_inst(
    .clk(clk),
    .reset(reset),
    .Instr(Instr[31:12]),
    .ALUFlags(ALUFlags),
    .RegSrc(RegSrc),
    .RegWrite(RegWrite),
    .ImmSrc(ImmSrc),
    .ALUSrc(ALUSrc),
    .ALUControl(ALUControl),
    .MemWrite(MemWrite),
    .MemtoReg(MemtoReg),
    .PCSrc(PCSrc),
    .DMSrc(DMSrc),
    .Shift(ShftOp),
    .Div(Division),
    .Mul(Multiplication),
    .Div_sel(DivMode),
    .Instrnew(NewInstr)
	);

    datapath datapath_inst(
        .clk(clk),
        .reset(reset),
        .RegSrc(RegSrc),
        .RegWrite(RegWrite),
        .ImmSrc(ImmSrc),
        .ALUSrc(ALUSrc),
        .ALUControl(ALUControl),
        .MemtoReg(MemtoReg),
        .PCSrc(PCSrc),
        .ALUFlags(ALUFlags),
        .PC(PC),
        .Instr(Instr),
        .ALUResult(ALUResult),
        .WriteData(WriteData),
        .ReadData(ReadData),
        .DMSrc(DMSrc),
    	.Shift(ShftOp),
    	.Div(Division),
    	.Mul(Multiplication),
    	.Div_sel(DivMode)
    	);
endmodule